library verilog;
use verilog.vl_types.all;
entity Control_Division_vlg_vec_tst is
end Control_Division_vlg_vec_tst;
