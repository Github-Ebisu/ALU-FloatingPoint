library verilog;
use verilog.vl_types.all;
entity Main_vlg_vec_tst is
end Main_vlg_vec_tst;
