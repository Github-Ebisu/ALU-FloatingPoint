library verilog;
use verilog.vl_types.all;
entity Mantissa_vlg_vec_tst is
end Mantissa_vlg_vec_tst;
