library verilog;
use verilog.vl_types.all;
entity FloatingPointMultiplication_vlg_vec_tst is
end FloatingPointMultiplication_vlg_vec_tst;
