library verilog;
use verilog.vl_types.all;
entity ALU_48bit_vlg_vec_tst is
end ALU_48bit_vlg_vec_tst;
