library verilog;
use verilog.vl_types.all;
entity Mantissa_Division_vlg_vec_tst is
end Mantissa_Division_vlg_vec_tst;
