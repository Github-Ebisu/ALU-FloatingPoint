library verilog;
use verilog.vl_types.all;
entity Mantissa_Division_vlg_sample_tst is
    port(
        A               : in     vl_logic_vector(22 downto 0);
        B               : in     vl_logic_vector(22 downto 0);
        CLK             : in     vl_logic;
        Start           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Mantissa_Division_vlg_sample_tst;
