library verilog;
use verilog.vl_types.all;
entity ALU_48bit_vlg_check_tst is
    port(
        Z               : in     vl_logic_vector(47 downto 0);
        sampler_rx      : in     vl_logic
    );
end ALU_48bit_vlg_check_tst;
